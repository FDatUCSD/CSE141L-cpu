`timescale 1ns / 1ps

module tb_ALU;

  // Inputs
  logic [2:0] OP;
  logic [7:0] R1, R2;

  // Outputs
  logic [7:0] OUT;
  logic [1:0] OVERFLOW;
  logic ZF;

  // Instantiate the ALU
  ALU uut (
    .OP(OP),
    .R1(R1),
    .R2(R2),
    .OUT(OUT),
    .OVERFLOW(OVERFLOW),
    .ZF(ZF)
  );

  // Task to display the result in binary
  task print_result(string op_name);
    $display("[%s] R1 = %08b, R2 = %08b => OUT = %08b, OVERFLOW = %02b, ZF = %b", 
             op_name, R1, R2, OUT, OVERFLOW, ZF);
  endtask

  initial begin
    $display("Starting ALU testbench...");

    // AND
    OP = 3'b000; R1 = 8'b10101010; R2 = 8'b11001100;
    #1; print_result("AND");

    // XOR
    OP = 3'b001; R1 = 8'b11110000; R2 = 8'b10101010;
    #1; print_result("XOR");

    // SHL (left shift R2 by R1 bits)
    OP = 3'b010; R1 = 3; R2 = 8'b00000001;
    #1; print_result("SHL");

    // SHR (right shift R2 by R1 bits)
    OP = 3'b011; R1 = 2; R2 = 8'b10000000;
    #1; print_result("SHR");

    // ADD (normal)
    OP = 3'b100; R1 = 8'd15; R2 = 8'd10;
    #1; print_result("ADD (normal)");

    // ADD (overflow)
    OP = 3'b100; R1 = 8'd255; R2 = 8'd255;
    #1; print_result("ADD (overflow)");

    // ADD (zero flag)
    OP = 3'b100; R1 = 8'd0; R2 = 8'd0;
    #1; print_result("ADD (ZF=1)");

    // Invalid OP (default case)
    OP = 3'b111; R1 = 8'hAA; R2 = 8'h55;
    #1; print_result("INVALID");

    $display("ALU testbench complete.");
  end

endmodule

